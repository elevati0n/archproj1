module controlunit ( output reg regdest, output reg jump, output reg branch, output reg memread,
                     output reg memtoreg, output reg memwrite, output reg alusrc, output reg regwrite,
                     output reg[1:0] aluop, input [5:0] opcode );
  // These cases and outputs are taken from figure 4.22, P&H 
  initial begin
      regdest = 0;
      alusrc = 0;
      memtoreg = 0;
      regwrite = 0;
      memread = 0;
      memwrite = 0;
      branch = 0;
      aluop = 2'b00;
      jump = 0;
  end 

                  
  always @ (opcode) begin
    {regdest, alusrc, memtoreg, regwrite, memread, memwrite, branch, jump, aluop}=10'b0000000000;
    case (opcode)
      6'b000000: begin // r-type, others are 0 by default
          regdest = 1;
          alusrc = 0;
          memtoreg = 0;
          regwrite = 1;
          memread = 0;
          memwrite = 0;
          branch = 0;
          aluop = 2'b10;
          jump = 0;
      end
      6'b100011: begin // lw
          regdest = 0;
          alusrc = 1;
          memtoreg = 0;
          regwrite = 1;
          memread = 1;
          memwrite = 0;
          branch = 0;
          aluop = 2'b00;
          jump = 0;
	end 
      6'b101011: begin // sw
        //regdest = x;
          alusrc = 1;
          memtoreg = 1;
          regwrite = 0;
          memread = 0;
          memwrite = 1;
          branch = 0;
          aluop = 2'b00;
          jump = 0;
       
      end
      6'b000100: begin // beq
        //regdest = x;
          alusrc = 0;
        //memtoreg = x;
          regwrite = 0;
          memread = 0;
          memwrite = 0;
          branch = 1;
          aluop = 2'b01;
          jump = 0;
      end
      6'b001000: begin // addi
          regdest = 0;
          alusrc = 1;
          memtoreg = 0;
          regwrite = 1;
          memread = 0;
          memwrite = 0;
          branch = 0;
          aluop = 2'b10;
          jump = 0;
      end
      6'b000010: begin // j
        jump = 1;
        // all else is don't-care
      end
     
    endcase
  end
endmodule
